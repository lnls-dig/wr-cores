library ieee;
use ieee.std_logic_1164.all;

package vfchd_i2cmux_pkg is

  component SfpIdReader is
    generic (
      g_SfpWbBaseAddress : natural := 0;
      g_WbAddrWidth      : natural := 32);
    port (
      Clk_ik       : in  std_logic;
      SfpPlugged_i : in  std_logic;
      SfpIdValid_o : out std_logic;
      SfpPN_b128   : out std_logic_vector(127 downto 0);
      WbCyc_o      : out std_logic;
      WbStb_o      : out std_logic;
      WbAddr_ob    : out std_logic_vector(g_WbAddrWidth-1 downto 0);
      WbData_ib8   : in  std_logic_vector(7 downto 0);
      WbAck_i      : in  std_logic);
  end component SfpIdReader;

  component I2cExpAndMuxMaster is
    generic (
      g_SclHalfPeriod : std_logic_vector(9 downto 0) := "0100000000");
    port (
      Clk_ik              : in    std_logic;
      Rst_irq             : in    std_logic;
      IoExpWrReq_i        : in    std_logic;
      IoExpWrOn_oq        : out   std_logic;
      IoExpRdReq_i        : in    std_logic;
      IoExpRdOn_oq        : out   std_logic;
      IoExpAddr_ib3       : in    std_logic_vector(2 downto 0);
      IoExpRegAddr_ib2    : in    std_logic_vector(1 downto 0);
      IoExpData_ib8       : in    std_logic_vector(7 downto 0);
      I2cSlaveWrReq_i     : in    std_logic;
      I2cSlaveWrOn_o      : out   std_logic;
      I2cSlaveRdReq_i     : in    std_logic;
      I2cSlaveRdOn_o      : out   std_logic;
      I2cMuxAddress_i     : in    std_logic;
      I2cMuxChannel_ib2   : in    std_logic_vector(1 downto 0);
      I2cSlaveAddr_ib7    : in    std_logic_vector(6 downto 0);
      I2cSlaveRegAddr_ib8 : in    std_logic_vector(7 downto 0);
      I2cSlaveByte_ib8    : in    std_logic_vector(7 downto 0);
      Busy_o              : out   std_logic;
      NewByteRead_op      : out   std_logic;
      ByteOut_ob8         : out   std_logic_vector(7 downto 0);
      AckError_op         : out   std_logic;
      Scl_ioz             : inout std_logic;
      Sda_ioz             : inout std_logic);
  end component I2cExpAndMuxMaster;

  component I2cExpAndMuxReqArbiter is
    port (
      Clk_ik                     : in  std_logic;
      Rst_irq                    : in  std_logic;
      IoExpWrReq_oq              : out std_logic;
      IoExpWrOn_i                : in  std_logic;
      IoExpRdReq_oq              : out std_logic;
      IoExpRdOn_i                : in  std_logic;
      IoExpAddr_oqb3             : out std_logic_vector(2 downto 0);
      IoExpRegAddr_oqb2          : out std_logic_vector(1 downto 0);
      IoExpData_oqb8             : out std_logic_vector(7 downto 0);
      I2cSlaveWrReq_oq           : out std_logic;
      I2cSlaveWrOn_i             : in  std_logic;
      I2cSlaveRdReq_oq           : out std_logic;
      I2cSlaveRdOn_i             : in  std_logic;
      I2cMuxAddress_oq           : out std_logic;
      I2cMuxChannel_oqb2         : out std_logic_vector(1 downto 0);
      I2cSlaveAddr_oqb7          : out std_logic_vector(6 downto 0);
      I2cSlaveRegAddr_oqb8       : out std_logic_vector(7 downto 0);
      I2cSlaveByte_oqb8          : out std_logic_vector(7 downto 0);
      MasterBusy_i               : in  std_logic;
      MasterNewByteRead_ip       : in  std_logic;
      MasterByteOut_ib8          : in  std_logic_vector(7 downto 0);
      MasterAckError_i           : in  std_logic;
      IoExpApp12Int_ian          : in  std_logic;
      IoExpApp34Int_ian          : in  std_logic;
      IoExpBstEthInt_ian         : in  std_logic;
      IoExpLosInt_ian            : in  std_logic;
      IoExpBlmInInt_ian          : in  std_logic;
      InitDone_oq                : out std_logic;
      VmeGa_onqb5                : out std_logic_vector(4 downto 0);
      VmeGaP_onq                 : out std_logic;
      Led_ib8                    : in  std_logic_vector(7 downto 0);
      StatusLed_ob8              : out std_logic_vector(7 downto 0);
      GpIo1A2B_i                 : in  std_logic;
      EnGpIo1Term_i              : in  std_logic;
      GpIo2A2B_i                 : in  std_logic;
      EnGpIo2Term_i              : in  std_logic;
      GpIo34A2B_i                : in  std_logic;
      EnGpIo3Term_i              : in  std_logic;
      EnGpIo4Term_i              : in  std_logic;
      StatusGpIo1A2B_oq          : out std_logic;
      StatusEnGpIo1Term_oq       : out std_logic;
      StatusGpIo2A2B_oq          : out std_logic;
      StatusEnGpIo2Term_oq       : out std_logic;
      StatusGpIo34A2B_oq         : out std_logic;
      StatusEnGpIo3Term_oq       : out std_logic;
      StatusEnGpIo4Term_oq       : out std_logic;
      BlmIn_oqb8                 : out std_logic_vector(7 downto 0);
      AppSfp1Present_oq          : out std_logic;
      AppSfp1Id_oq16             : out std_logic_vector(15 downto 0);
      AppSfp1TxFault_oq          : out std_logic;
      AppSfp1Los_oq              : out std_logic;
      AppSfp1TxDisable_i         : in  std_logic;
      AppSfp1RateSelect_i        : in  std_logic;
      StatusAppSfp1TxDisable_oq  : out std_logic;
      StatusAppSfp1RateSelect_oq : out std_logic;
      AppSfp2Present_oq          : out std_logic;
      AppSfp2Id_oq16             : out std_logic_vector(15 downto 0);
      AppSfp2TxFault_oq          : out std_logic;
      AppSfp2Los_oq              : out std_logic;
      AppSfp2TxDisable_i         : in  std_logic;
      AppSfp2RateSelect_i        : in  std_logic;
      StatusAppSfp2TxDisable_oq  : out std_logic;
      StatusAppSfp2RateSelect_oq : out std_logic;
      AppSfp3Present_oq          : out std_logic;
      AppSfp3Id_oq16             : out std_logic_vector(15 downto 0);
      AppSfp3TxFault_oq          : out std_logic;
      AppSfp3Los_oq              : out std_logic;
      AppSfp3TxDisable_i         : in  std_logic;
      AppSfp3RateSelect_i        : in  std_logic;
      StatusAppSfp3TxDisable_oq  : out std_logic;
      StatusAppSfp3RateSelect_oq : out std_logic;
      AppSfp4Present_oq          : out std_logic;
      AppSfp4Id_oq16             : out std_logic_vector(15 downto 0);
      AppSfp4TxFault_oq          : out std_logic;
      AppSfp4Los_oq              : out std_logic;
      AppSfp4TxDisable_i         : in  std_logic;
      AppSfp4RateSelect_i        : in  std_logic;
      StatusAppSfp4TxDisable_oq  : out std_logic;
      StatusAppSfp4RateSelect_oq : out std_logic;
      BstSfpPresent_oq           : out std_logic;
      BstSfpId_oq16              : out std_logic_vector(15 downto 0);
      BstSfpTxFault_oq           : out std_logic;
      BstSfpLos_oq               : out std_logic;
      BstSfpTxDisable_i          : in  std_logic;
      BstSfpRateSelect_i         : in  std_logic;
      StatusBstSfpTxDisable_oq   : out std_logic;
      StatusBstSfpRateSelect_oq  : out std_logic;
      EthSfpPresent_oq           : out std_logic;
      EthSfpId_oq16              : out std_logic_vector(15 downto 0);
      EthSfpTxFault_oq           : out std_logic;
      EthSfpLos_oq               : out std_logic;
      EthSfpTxDisable_i          : in  std_logic;
      EthSfpRateSelect_i         : in  std_logic;
      StatusEthSfpTxDisable_oq   : out std_logic;
      StatusEthSfpRateSelect_oq  : out std_logic;
      CdrLos_oq                  : out std_logic;
      CdrLol_oq                  : out std_logic;
      I2cWbCyc_i                 : in  std_logic;
      I2cWbStb_i                 : in  std_logic;
      I2cWbWe_i                  : in  std_logic;
      I2cWbAdr_ib12              : in  std_logic_vector(11 downto 0);
      I2cWbDat_ib8               : in  std_logic_vector(7 downto 0);
      I2cWbDat_ob8               : out std_logic_vector(7 downto 0);
      I2cWbAck_o                 : out std_logic;
      WbCyc_i                    : in  std_logic;
      WbStb_i                    : in  std_logic;
      WbWe_i                     : in  std_logic;
      WbDat_ib32                 : in  std_logic_vector(31 downto 0);
      WbDat_oqb32                : out std_logic_vector(31 downto 0);
      WbAck_oa                   : out std_logic);
  end component I2cExpAndMuxReqArbiter;

end vfchd_i2cmux_pkg;
