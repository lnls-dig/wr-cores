`define ADDR_WRC_DIAGS_CTRL            7'h0
`define WRC_DIAGS_CTRL_DATA_VALID_OFFSET 0
`define WRC_DIAGS_CTRL_DATA_VALID 32'h00000001
`define WRC_DIAGS_CTRL_DATA_SNAPSHOT_OFFSET 8
`define WRC_DIAGS_CTRL_DATA_SNAPSHOT 32'h00000100
`define ADDR_WRC_DIAGS_WDIAG_SSTAT     7'h4
`define WRC_DIAGS_WDIAG_SSTAT_WR_MODE_OFFSET 0
`define WRC_DIAGS_WDIAG_SSTAT_WR_MODE 32'h00000001
`define WRC_DIAGS_WDIAG_SSTAT_SERVOSTATE_OFFSET 8
`define WRC_DIAGS_WDIAG_SSTAT_SERVOSTATE 32'h00000f00
`define ADDR_WRC_DIAGS_WDIAG_PSTAT     7'h8
`define WRC_DIAGS_WDIAG_PSTAT_LINK_OFFSET 0
`define WRC_DIAGS_WDIAG_PSTAT_LINK 32'h00000001
`define WRC_DIAGS_WDIAG_PSTAT_LOCKED_OFFSET 1
`define WRC_DIAGS_WDIAG_PSTAT_LOCKED 32'h00000002
`define ADDR_WRC_DIAGS_WDIAG_PTPSTAT   7'hc
`define WRC_DIAGS_WDIAG_PTPSTAT_PTPSTATE_OFFSET 0
`define WRC_DIAGS_WDIAG_PTPSTAT_PTPSTATE 32'h000000ff
`define ADDR_WRC_DIAGS_WDIAG_ASTAT     7'h10
`define WRC_DIAGS_WDIAG_ASTAT_AUX_OFFSET 0
`define WRC_DIAGS_WDIAG_ASTAT_AUX 32'h000000ff
`define ADDR_WRC_DIAGS_WDIAG_TXFCNT    7'h14
`define ADDR_WRC_DIAGS_WDIAG_RXFCNT    7'h18
`define ADDR_WRC_DIAGS_WDIAG_SEC_MSB   7'h1c
`define ADDR_WRC_DIAGS_WDIAG_SEC_LSB   7'h20
`define ADDR_WRC_DIAGS_WDIAG_NS        7'h24
`define ADDR_WRC_DIAGS_WDIAG_MU_MSB    7'h28
`define ADDR_WRC_DIAGS_WDIAG_MU_LSB    7'h2c
`define ADDR_WRC_DIAGS_WDIAG_DMS_MSB   7'h30
`define ADDR_WRC_DIAGS_WDIAG_DMS_LSB   7'h34
`define ADDR_WRC_DIAGS_WDIAG_ASYM      7'h38
`define ADDR_WRC_DIAGS_WDIAG_CKO       7'h3c
`define ADDR_WRC_DIAGS_WDIAG_SETP      7'h40
`define ADDR_WRC_DIAGS_WDIAG_UCNT      7'h44
`define ADDR_WRC_DIAGS_WDIAG_TEMP      7'h48
